`include "CPU_define.vh"

module CPU_bank_reg
(
    input wire clock,
    input wire reset,
    
    CPU_bank_reg_if.slave bank_reg_if
);

integer i;
reg [`REG_WIDTH-1:0] reg_file [`NUM_REGS];

always @(posedge clock) begin
    if (reset) begin 
        for (i=0; i<`NUM_REGS; i=i+1) reg_file[i] <= 0;
    end else begin
        bank_reg_if.read_data_a <= reg_file[bank_reg_if.read_reg_a];
        bank_reg_if.read_data_b <= reg_file[bank_reg_if.read_reg_b];
        if (bank_reg_if.write_enable) reg_file[bank_reg_if.write_reg] <= bank_reg_if.write_data;
    end
end

endmodule
